library verilog;
use verilog.vl_types.all;
entity tb_LFSR is
end tb_LFSR;
